module goodbye_world ;

initial begin
  $display ("Goodbye World");
   #10  $finish;
end

endmodule
